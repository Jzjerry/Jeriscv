module TopLevel();
    
endmodule